library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

library work;
use work.common.all;

entity imem is
    port(
        addr : in std_logic_vector(6 downto 0);
        dout : out word);
end imem;

architecture behavioral of imem is
type rom_arr is array(0 to 127) of word;
--00010224 T main
constant mem:rom_arr:=
    (
    --tausseed
   x"00a02823", --  		sw	a0,16(zero)
   x"00002A23", --  		sw	zero,20(zero)
   x"00002C23", --  		sw	zero,24(zero)
   x"00008067", --  67800000 		ret
   x"00000013", --  13000000                nop
   --taus
   x"01002783", --  		lw	a5,16(zero)
   x"00000013", --       13000000                nop
   x"00D79513", -- 1395D700 		slli	a0,a5,13
   x"00F54533", -- 3345F500 		xor	a0,a0,a5
   x"01355513", -- 13553501 		srli	a0,a0,19
   x"00C79793", -- 9397C700 		slli	a5,a5,12
   x"FFFFE6B7", -- B7E6FFFF 		li	a3,-8192
   x"00D7F7B3", -- B3F7D700 		and	a5,a5,a3
   x"00F54533", -- 3345F500 		xor	a0,a0,a5
   x"00000013", --       13000000                nop
   x"00a02823", --  		sw	a0,16(zero)
   x"01402783", --  		lw	a5,20(zero)
   x"00000013", --       13000000                nop
   x"00279713", -- 13972700 		slli	a4,a5,2
   x"00F74733", -- 3347F700 		xor	a4,a4,a5
   x"01975713", -- 13579701 		srli	a4,a4,25
   x"00479793", -- 93974700 		slli	a5,a5,4
   x"F807F793", -- 93F707F8 		andi	a5,a5,-128
   x"00F74733", -- 3347F700 		xor	a4,a4,a5
   x"00000013", --       13000000                nop
   x"00E02A23", --  		sw	a4,20(zero)
   x"01802783", --  		lw	a5,24(zero)
   x"00000013", --       13000000                nop
   x"00379693", -- 93963700 		slli	a3,a5,3
   x"00F6C6B3", -- B3C6F600 		xor	a3,a3,a5
   x"00B6D693", -- 93D6B600 		srli	a3,a3,11
   x"01179793", -- 93971701 		slli	a5,a5,17
   x"FFE005B7", -- B705E0FF 		li	a1,-2097152
   x"00B7F7B3", -- B3F7B700 		and	a5,a5,a1
   x"00D7C7B3", -- B3C7D700 		xor	a5,a5,a3
   x"00000013", --       13000000                nop
   x"00F02C23", --  		sw	a5,24(zero)
   x"00E54533", -- 3345E500 		xor	a0,a0,a4
   x"00F54533", -- 3345F500 		xor	a0,a0,a5
   x"00008067", --67800000 		ret
   x"00000013", --       13000000                nop
   --main
   x"FF010113", -- 130101FF 		addi	sp,sp,-16
   x"00000013", --       13000000                nop
   x"00112623", -- 23261100 		sw	ra,12(sp)
   x"00812423", -- 23248100 		sw	s0,8(sp)
   x"00912223", -- 23229100 		sw	s1,4(sp)
   x"01212023", -- 23202101 		sw	s2,0(sp)
   x"1C9F0537", -- 3765BC00 		lui a0, 0x1c9f0
   x"79250513", -- 1305E514 		addi	a0,a0,1938
   x"F39FF0EF", -- 97000000 		jal   pc - 0xa0 call tausseed
   x"00000013", --       13000000                nop
   x"00000413", -- 13040000 		li	s0,0
   x"01400493", -- 93044001 		li	s1,20
   --L4 loop starts here
   x"F3DFF0EF", --  		jal     pc - 0xa0  call	taus
   x"00000013", --       13000000                nop
   x"00050613", -- 13060500 		mv	a2,a0
   x"00040593", -- 93050400 		mv	a1,s0
   x"00140413", -- 13041400 		addi	s0,s0,1
   x"00000013", --       13000000                nop
   x"FE9412E3", --  		bne	s0,s1,.L4
   x"00000013", --       13000000                nop
   x"00000513", -- 13050000 		li	a0,0
   x"00C12083", -- 8320C100 		lw	ra,12(sp)
   x"00812403", -- 03248100 		lw	s0,8(sp)
   x"00412483", -- 83244100 		lw	s1,4(sp)
   x"00012903", -- 03290100 		lw	s2,0(sp)
   x"01010113", -- 13010101 		addi	sp,sp,16
   x"00008067",
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013", --       13000000                nop
   x"00000013"); -- ret


begin
	dout<=mem(conv_integer(addr));
end behavioral;
